LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY KALKULATOR IS
GENERIC ( N : NATURAL := 2);
PORT(	
	 CLK        : IN 		STD_LOGIC;
    A          : INOUT 	INTEGER RANGE 0 TO 100;
    B        	: INOUT 	INTEGER RANGE 0 TO 100;
    SUM       	: OUT 	INTEGER RANGE 0 TO 999999;
	 SUM2    	: OUT 	INTEGER RANGE 0 TO 999999;
    MODE       : IN 		INTEGER RANGE 0 TO 1;
	 SEL1  		: IN 		INTEGER RANGE 0 TO 7;
	 SEL2  		: IN 		INTEGER RANGE 0 TO 8);
END KALKULATOR;

ARCHITECTURE HASIL OF KALKULATOR IS
SIGNAL TEMPADD        : INTEGER;
SIGNAL TEMPSUB        : INTEGER;
SIGNAL TEMPMUL        : INTEGER;
SIGNAL TEMPDIV        : INTEGER;
SIGNAL TEMPROOT       : INTEGER;
SIGNAL TEMPROOT2      : INTEGER:=11;
SIGNAL TEMPPOW        : INTEGER;
SIGNAL MS_TO_KMH   	 : INTEGER;
SIGNAL C_TO_K    		 : INTEGER;
SIGNAL C_TO_R   		 : INTEGER;
SIGNAL C_TO_F    		 : INTEGER;
SIGNAL H_TO_S	    	 : INTEGER;
SIGNAL DISTANCE		 : INTEGER;
SIGNAL DEBIT			 : INTEGER;
SIGNAL VOLT				 : INTEGER;
SIGNAL PECAHAN_BULAT	 : INTEGER;
SIGNAL PECAHAN_KOMA	 : INTEGER;
SIGNAL SQRTROOT		 : INTEGER:=10;

BEGIN
PROCESS (CLK, MODE, SEL1, SEL2)
BEGIN 
	IF(RISING_EDGE(CLK) AND MODE = 0) THEN 
		CASE SEL1 IS  
			WHEN 0 => A	<=0; B <= 0;SUM <= 0;SUM2 <= 0;TEMPADD <= 0;TEMPSUB <= 0;TEMPMUL <= 0;TEMPDIV <= 0;TEMPROOT <= 0;
						 TEMPPOW <= 0;PECAHAN_BULAT <= 0;PECAHAN_KOMA <= 0;PECAHAN_KOMA <= 0;SQRTROOT	<= 0;TEMPROOT2 <= 11;
						 SQRTROOT	<= 10;
			WHEN 1 => TEMPADD <= A + B; SUM <= TEMPADD;
			WHEN 2 => TEMPSUB <= A - B; SUM <= TEMPSUB;
			WHEN 3 => TEMPMUL <= A * B; SUM <= TEMPMUL;
			WHEN 4 => TEMPDIV <= A / B; SUM <= TEMPDIV;
			WHEN 5 => PECAHAN_BULAT  <= A / B;	
						 PECAHAN_KOMA   <= ((A - (B*PECAHAN_BULAT)) * 10) / B;
						 SUM 				 <= PECAHAN_BULAT;--STORE PECAHAN ANGKA BULAT (...,00)
						 SUM2 			 <= PECAHAN_KOMA;	--STORE PECAHAN ANGKA DIBELAKANG KOMA (1,000)
			WHEN 6 => TEMPPOW <= A ** N; SUM <= TEMPPOW;
			WHEN 7 => FOR I IN 1 TO 10 LOOP		--AKAR DARI NILAI A
						 TEMPROOT <= SQRTROOT**N;
							IF TEMPROOT = A THEN	SUM<= TEMPROOT2;
							EXIT;
							ELSIF TEMPROOT < A THEN	SUM<= TEMPROOT2;		
							EXIT;
							END IF;
						 TEMPROOT2<=TEMPROOT2-1;
						 SQRTROOT<=SQRTROOT-1;
						 END LOOP;
						 FOR I IN 1 TO 10 LOOP		--AKAR DARI NILAI B
						 TEMPROOT <= SQRTROOT**N;
							IF TEMPROOT = B THEN	SUM2<= TEMPROOT2;
							EXIT;
							ELSIF TEMPROOT < B THEN	SUM2<= TEMPROOT2;		
							EXIT;
							END IF;
						 TEMPROOT2<=TEMPROOT2-1;
						 SQRTROOT<=SQRTROOT-1;
						 END LOOP;
		END CASE;
	ELSIF(RISING_EDGE(CLK) AND MODE = 1) THEN 
		CASE SEL2 IS
			WHEN 0 => A	<= 0;B <= 0;SUM <= 0;MS_TO_KMH <= 0; C_TO_K <= 0; C_TO_R<= 0;C_TO_F <= 0;H_TO_S	<= 0;DISTANCE <= 0;
						 DEBIT <= 0; VOLT <= 0;	
			WHEN 1 => MS_TO_KMH 	<= ((A *18)/5); SUM <= MS_TO_KMH;
			WHEN 2 => C_TO_K 		<= (A + 273); SUM <= C_TO_K;
			WHEN 3 => C_TO_R 		<= ((A*4)/5); SUM <= C_TO_R;
			WHEN 4 => C_TO_F  	<= (((A *9)/5)+32); SUM <= C_TO_F;
			WHEN 5 => H_TO_S  	<= (A *3600); SUM <= H_TO_S;
			WHEN 6 => DISTANCE  	<= (A *B);--SPEED* TIME 
						 SUM 			<= DISTANCE;--A=SPEED, B=TIME
			WHEN 7 => DEBIT  		<= (A/B); --VOLUME/TIME
						 SUM 			<= DEBIT;
			WHEN 8 => VOLT 		<= (A*B);--VOLT= I * R
						 SUM 			<= VOLT;
		END CASE;
	END IF;
END PROCESS;
END HASIL;